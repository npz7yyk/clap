module csr
(
    input clk,rstn
);

endmodule
