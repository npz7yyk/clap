// -*- Verilog -*-

`ifdef VERILATOR
`define CLAP_CONFIG_DIFFTEST
`define CLAP_CONFIG_BR_PROFILE
`define CLAP_CONFIG_INST_PROFILE
`endif
