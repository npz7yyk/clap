// -*- Verilog -*-

`ifdef VERILATOR
`define CLAP_CONFIG_DIFFTEST
`define CLAP_CONFIG_BR_PROFILE
`define CLAP_CONFIG_INST_PROFILE
`define CLAP_CONFIG_AXI_PROFILE
`define CLAP_CONFIG_LD_ST_PROFILE
`endif
