`timescale 1ns / 1ps

module TagV_memory(
    input clk,
    input [31:0] r_addr,
    input [31:0] w_addr,
    input [3:0] we,
    output [3:0] hit,
    output cache_hit
    );
    wire [5:0] index;
    wire [19:0] tag;
    wire [19:0] tag_0, tag_1, tag_2, tag_3;
    wire vld_0, vld_1, vld_2, vld_3;

    assign index = r_addr[11:6];
    assign tag = r_addr[31:12];

    assign hit[0] = (tag == tag_0) && vld_0;
    assign hit[1] = (tag == tag_1) && vld_1;
    assign hit[2] = (tag == tag_2) && vld_2;
    assign hit[3] = (tag == tag_3) && vld_3;

    assign cache_hit = |hit;
    TagV way0_TagV(
        .addra  (index),
        .clka   (clk),
        .dina   ({1'b1, w_addr[31:12]}),
        .wea    (we[0]),
        .addrb  (index),
        .clkb   (clk),
        .doutb  ({vld_0, tag_0})
    );
    TagV way1_TagV(
        .addra  (index),
        .clka   (clk),
        .dina   ({1'b1, w_addr[31:12]}),
        .wea    (we[1]),
        .addrb  (index),
        .clkb   (clk),
        .doutb  ({vld_1, tag_1})
    );
    TagV way2_TagV(
        .addra  (index),
        .clka   (clk),
        .dina   ({1'b1, w_addr[31:12]}),
        .wea    (we[2]),
        .addrb  (index),
        .clkb   (clk),
        .doutb  ({vld_2, tag_2})
    );
    TagV way3_TagV(
        .addra  (index),
        .clka   (clk),
        .dina   ({1'b1, w_addr[31:12]}),
        .wea    (we[3]),
        .addrb  (index),
        .clkb   (clk),
        .doutb  ({vld_3, tag_3})
    );

endmodule
